LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

ENTITY controller IS
	PORT (
		IR : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		SW : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
		S : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		SEL : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		W1, W2, W3, T3, C, Z, CLR : IN STD_LOGIC;
		LIR, PCINC, ARINC, PCADD, M, CIN, ABUS, DRW, MEMW, LDZ, LDC, LAR, LONG, SHORT, MBUS, SBUS, LPC, SELCTL, STOP : OUT STD_LOGIC
	);
END controller;

ARCHITECTURE behaviour OF controller IS
	-- Temp Variable Definition
	SIGNAL ST0 : STD_LOGIC; -- indicate next stage
	SIGNAL SST0 : STD_LOGIC; -- indicate change of ST0
BEGIN
	-- Behaviour of Controller
	-- CLR & T3 occurs
	PROCESS (CLR, T3)
	BEGIN
		IF (T3'EVENT AND T3 = '0' AND SST0 = '1') THEN -- descending edge of T3
			ST0 <= '1'; -- Indicate Stage 2
		END IF;

		IF (CLR = '0') THEN
			ST0 <= '0'; -- Default ST0
		END IF;
	END PROCESS;

	-- Other signals change
	PROCESS (SW, W1, W2, W3, IR, C, Z, ST0)
	BEGIN
		-- Initialize all output signals
		LIR <= '0';
		PCINC <= '0';
		ARINC <= '0';
		PCADD <= '0';
		M <= '0';
		S <= "0000";
		SEL <= "0000";
		CIN <= '0';
		ABUS <= '0';
		SBUS <= '0';
		DRW <= '0';
		MEMW <= '0';
		LDZ <= '0';
		LDC <= '0';
		LAR <= '0';
		LONG <= '0';
		SHORT <= '0';
		MBUS <= '0';
		LPC <= '0';
		SELCTL <= '0';
		STOP <= '0';

		SST0 <= '0'; -- Default SST0

		CASE SW IS
			WHEN "001" => -- Write into Mem
				SBUS <= W1;
				LAR <= (NOT ST0) AND W1;
				STOP <= W1;
				SST0 <= (NOT ST0) AND W1;
				SHORT <= W1;
				SELCTL <= W1;
				MEMW <= (ST0) AND W1;
				ARINC <= (ST0) AND W1;
			WHEN "010" => -- Read from mem
				SBUS <= (NOT ST0) AND W1;
				LAR <= (NOT ST0) AND W1;
				STOP <= W1;
				SST0 <= (NOT ST0) AND W1;
				SHORT <= W1;
				SELCTL <= W1;
				MBUS <= (ST0) AND W1;
				ARINC <= (ST0) AND W1;
			WHEN "011" => -- Read from reg
				SEL <= ((NOT W1) AND W2) & '0' & ((NOT W1) AND W2) & '1';
				SELCTL <= W1 OR W2;
				STOP <= W1 OR W2;
			WHEN "100" => -- Write into reg
				SBUS <= W1 or W2;
				SEL <= ST0 & W2 & (((NOT ST0) AND W1) OR (ST0 AND W2)) & W1;
				DRW <= W1 OR W2;
				STOP <= W1 OR W2;
				SELCTL <= W1 OR W2;
				SST0 <= (NOT ST0) AND W2;
			WHEN "000" => -- Instruction Fetching
				IF ST0 = '0' THEN -- Stage 1: Read from user input, write into PC
					SST0 <= W1; -- Indicate ST0='1' next round
					LPC <= W1;
					SHORT <= W1; -- Restart from W1 next round
					SBUS <= W1; -- Read from keyboard
					-- STOP <= '1'; -- Try stop
				ELSE -- Stage 2: Read from given addr
					CASE IR IS
						WHEN "0000"=> -- Initial State
							LIR <= W1;
							PCINC <= W1;
							SHORT <= W1; -- Restart from W1 next round
						WHEN "0001" => -- ADD
							S <= "1001";
							CIN <= W1; -- Perform A + B, A chosen by IR[3:2], B chosen by IR[1:0]
							ABUS <= W1;
							DRW <= W1; -- Write result into register(selected by IR[3:2])
							LDZ <= W1; -- Save the zero generated by the operation to the Z flag register on the rising edge of T3
							LDC <= W1; -- Save the carry generated by the operation to the C flag register on the rising edge of T3

							LIR <= W1;
							PCINC <= W1; -- Fetch next instruction in advance
							SHORT <= W1; -- Restart from W1 next round
						WHEN "0010" => -- SUB
							S <= "0110"; -- Perform A - B, A chosen by IR[3:2], B chosen by IR[1:0]
							ABUS <= W1;
							DRW <= W1; -- Write result into register(selected by IR[3:2])
							LDZ <= W1; -- Save the zero generated by the operation to the Z flag register on the rising edge of T3
							LDC <= W1; -- Save the carry generated by the operation to the C flag register on the rising edge of T3

							LIR <= W1;
							PCINC <= W1; -- Fetch next instruction in advance
							SHORT <= W1; -- Restart from W1 next round
						WHEN "0011" => -- AND
							M <= W1;
							S <= "1011"; -- Perform A AND B, A chosen by IR[3:2], B chosen by IR[1:0]
							ABUS <= W1;
							DRW <= W1; -- Write result into register(selected by IR[3:2])
							LDZ <= W1; -- Save the zero generated by the operation to the Z flag register on the rising edge of T3

							LIR <= W1;
							PCINC <= W1; -- Fetch next instruction in advance
							SHORT <= W1; -- Restart from W1 next round
						WHEN "0100" => --INC
							S <= "0000"; -- Perform A + 1, A chosen by IR[3:2], B = 1
							ABUS <= W1;
							DRW <= W1; -- Write result into register(selected by IR[3:2])
							LDZ <= W1;
							LDC <= W1;

							LIR <= W1;
							PCINC <= W1; -- Fetch next instruction in advance
							SHORT <= W1; -- Restart from W1 next round
						WHEN "0101" => -- LD
							-- Step 1: Write B port(selected by IR[1:0]) into AR
							M <= W1; 
							S <= "1010";
							ABUS <= W1;
							LAR <= W1;
							LONG <= W1;

							-- Step 2: Write MEM[AR] into register(selected by IR[3:2])
							DRW <= W2;
							MBUS <= W2;
							
							LIR <= W2;
							PCINC <= W2; -- Fetch next instruction in advance
						WHEN "0110" => -- ST
							-- Step 1: Write A port(IR[3:2]) into AR
							M <= W1 OR W2;
							S <= '1' & (W1 AND (NOT W2)) & '1' & (W1 AND (NOT W2));
							ABUS <= W1 OR W2;
							LAR <= W1;
							LONG <= W1;

							-- Equivalent code to IF code segment above
							-- IF statement will introduce a multiplexer, which is less efficient
							MEMW <= W2;
												
							LIR <= W2;
							PCINC <= W2; -- Fetch next instruction in advance
						WHEN "0111" => -- JC
							-- Equivalent code to IF code segment above
							-- IF statement will introduce a multiplexer, which is less efficient
							PCADD <= C AND W1; -- Jump instruction, can not directly use pipeline
							
							SHORT <= NOT C AND W1; -- Restart from W1 next round if there is no JUMP CAUSED BY JC
							LIR <= ((NOT C) AND W1) OR W2;
							PCINC <= ((NOT C) AND W1) OR W2; 
						WHEN "1000" => -- JZ
							-- Equivalent code to IF code segment above
							-- IF statement will introduce a multiplexer, which is less efficient
							PCADD <= Z AND W1;
							
							SHORT <= NOT Z AND W1; -- Restart from W1 next round if there is no JUMP CAUSED BY JZ
							LIR <= ((NOT Z) AND W1) OR W2;
							PCINC <= ((NOT Z) AND W1) OR W2; 
						WHEN "1001" => --JMP
							M <= W1;
							S <= "1111"; -- Select A port(chosen by IR[3:2])
							ABUS <= W1;
							LPC <= W1; -- Write A port into PC 

							LIR <= W2;
							PCINC <= W2; 
						WHEN "1110" => --STP
							STOP <= W1;

						-- Added Instructions
						WHEN "1010" => --OUT
							M <= W1;
							S <= "1010"; -- Select B port(chosen by IR[1:0])
							ABUS <= W1; -- Deliver B port to DBUS

							LIR <= W1;
							PCINC <= W1; -- Fetch next instruction in advance
							SHORT <= W1; -- Restart from W1 next round
						when "1011" => -- XOR
							S <= '0110'; -- Perform A XOR B, A chosen by IR[3:2], B chosen by IR[1:0]
							M <= W1;
							ABUS <= W1;
							DRW <= W1;
							LDZ <= W1;

							LIR <= W1;
							PCINC <= W1; -- Fetch next instruction in advance
							SHORT <= W1; -- Restart from W1 next round
						when "1100" => -- OR
							S <= '1110' -- Perform A OR B, A chosen by IR[3:2], B chosen by IR[1:0]
							M <= W1;
							ABUS <= W1; 
							DRW <= W1;
							LDZ <= W1;

							LIR <= W1; 
							PCINC <= W1; -- Fetch next instruction in advance
							SHORT <= W1; -- Restart from W1 next round
						when "1101" =>  -- NOT
							S <= '0000'; -- Perform NOT A, A chosen by IR[3:2]
							M <= W1;
							ABUS <= W1;
							DRW <= W1;
							LDZ <= W1;

							LIR <= W1;
							PCINC <= W1; -- Fetch next instruction in advance
							SHORT <= W1; -- Restart from W1 next round
						WHEN OTHERS =>
							NULL;
					END CASE;
				END IF;
			WHEN OTHERS =>
				NULL;
		END CASE;
	END PROCESS;
END behaviour;